// Code your testbench here
// or browse Examples
`include "pipe_pkg.sv"
`include "top.sv"