module pipe{ clk, 
rst_n,
i_cf,
i_en,
i_data0,i_data1,
o_data0,
o_data1
};

























endmodule
