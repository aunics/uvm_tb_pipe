
package pipe_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "transfer.sv" 
`include "pipe_driver.sv" 
`include "pipe_monitor.sv" 
`include "pipe_sequencer.sv" 
`include "pipe_scoreboard.sv" 
`include "pipe_agent.sv"
`include "pipe_env.sv" 
`include "dut_env.sv" 
`include "pipe_seqlib.sv"
`include "pipe_test.sv"
endpackage // pipe_pkg